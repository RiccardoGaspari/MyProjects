
.model NMOS NMOS(LEVEL=1, VTO=0.71, KP=182e-6, GAMMA=0.01, LAMBDA=0.01, PHI=0.6, tox=9.6e-9, cj=350e-6, cjsw=120e-12, pb=0.8, mj=0.33, mjsw=0.33, cgso=0.046e-9, cgdo=0.046e-9 )
.model PMOS PMOS(LEVEL=1, VTO=-0.901, KP=41.5e-6, GAMMA=0.01, LAMBDA=0.01, PHI=0.6, tox=9.6e-9, cj=350e-6, cjsw=120e-12, pb=0.8, mj=0.33, mjsw=0.33, cgso=0.046e-9, cgdo=0.046e-9 )

* Mx Drain Gate Source Bulk L= W=


.SUBCKT OPAMPF2022 3 2 8

* coppia differenziale
M1 4 2 1 10 NMOS L=1u W=0.84u
M2 6 3 1 10 NMOS L=1u W=0.84u

* specchio di corrente
M3 4 4 5 5 PMOS L=1u W=1u
M4 6 4 5 5 PMOS L=1u W=1u

* stadio di uscita
M6 8 6 5 5 PMOS L=17.7n W=0.27u
M7 8 9 10 10 NMOS L=1u W=2.9u

* circuito di polarizzazione
M5 1 9 10 10 NMOS L=1u W=0.39u
M8 9 9 10 10 NMOS L=1u W=50n
M14 11 9 13 10 NMOS L=1u W=70n

M10 9 11 14 5 PMOS L=1u W=0.27u
M11 14 12 5 5 PMOS L=1u W=0.27u
M13 12 12 5 5 PMOS L=1u W=0.27u
M12 11 11 12 5 PMOS L=1u W=0.27u

Rb 13 10 100k

* tensioni di alimentazione
Vdd 5 0 2.5V
Vss 0 10 2.5V


* compensazione
M9 7 11 6 5 PMOS L=1u W=2.1u
Cc 8 7 0.776p

CL 8 0 5p

*.OP

.ENDS OPAMPF2022


*
